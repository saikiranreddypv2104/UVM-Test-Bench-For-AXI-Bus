`include "uvm_macros.svh"
import uvm_pkg::*;
`include "transaction.sv"
`include "slave_transaction.sv"
`include "slave_driver.sv"
`include "slave_monitor.sv"
`include "slave_agent.sv"
`include "sequence.sv"
`include "driver.sv"
`include "monitor.sv"
`include "scoreboard.sv"
`include "agent.sv"
`include "env.sv"
`include "test.sv"